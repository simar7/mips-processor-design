module decode(clock, insn, pc);

endmodule
