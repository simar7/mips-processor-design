module decode(clock, insn, pc);

// Input ports
input clock;
input [31:0] insn;
input [31:0] pc;

// Registers
reg [31:0] pc_reg;

always @(posedge clock)
begin : DECODE

	

endmodule
